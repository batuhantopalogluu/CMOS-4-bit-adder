* CMOS NAND2
* BATUHAN TOPALOĞLU 2019 
* SPICE3 file created from nand2.ext - technology: scmos

.option scale=0.12u


M1000 out a vdd w_n8_8# pmos w=20 l=2
+  ad=120 pd=52 as=200 ps=100
M1001 vdd b out w_n8_8# pmos w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_5_n6# a gnd gnd nmos w=8 l=2
+  ad=48 pd=28 as=40 ps=26
M1003 out b a_5_n6# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0

C0 b w_n8_8# 0.09fF
C1 gnd out 0.04fF
C2 a w_n8_8# 0.09fF
C3 out w_n8_8# 0.06fF
C4 out vdd 0.49fF
C5 vdd w_n8_8# 0.21fF
C6 b a 0.07fF
C7 out b 0.02fF
C8 gnd gnd 0.20fF
C9 out gnd 0.07fF
C10 vdd gnd 0.05fF
C11 b Gnd 0.09fF
C12 a Gnd 0.09fF
C13 w_n8_8# gnd 0.99fF

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node  OptionT1  V1   T2  V2   T3   V3   T4  V4    T5   V5  T6   V6   T7   V7  T8  V8  T9   V9 
*----- ----- ----- ------ --  --   --  --  ---- --    --  --   ---- ---  --- ---  ---- ---
Vin     a     GND    PWL( 0   0    4N  0   4.1N  2.5  8N  2.5  8.1N  0  12N   0  12.1N  2.5 16N 2.5 16.1N 0) 
Vin2    b     GND    PWL( 0   0    4N  0   4.1N   0   8N   0   8.1N 2.5 12N  2.5 12.1N  2.5 16N 2.5 16.1N 0) 

*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd    gnd     DC=2.5

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  16.1N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
