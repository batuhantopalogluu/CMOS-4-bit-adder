magic
tech scmos
timestamp 1578055772
<< nwell >>
rect -8 8 16 42
<< ntransistor >>
rect 3 -6 5 2
<< ptransistor >>
rect 3 14 5 34
<< ndiffusion >>
rect 2 -6 3 2
rect 5 -6 6 2
<< pdiffusion >>
rect 2 14 3 34
rect 5 14 6 34
<< ndcontact >>
rect -2 -6 2 2
rect 6 -6 10 2
<< pdcontact >>
rect -2 14 2 34
rect 6 14 10 34
<< polysilicon >>
rect 3 34 5 37
rect 3 2 5 14
rect 3 -9 5 -6
<< polycontact >>
rect -8 6 3 10
<< metal1 >>
rect -8 38 16 42
rect -2 34 2 38
rect 6 10 10 14
rect 6 6 16 10
rect 6 2 10 6
rect -2 -10 2 -6
rect -8 -14 16 -10
<< labels >>
rlabel metal1 0 39 0 39 5 vdd
rlabel polycontact 0 8 0 8 1 a
rlabel metal1 12 8 12 8 7 y
rlabel metal1 4 -12 4 -12 1 gnd
<< end >>
