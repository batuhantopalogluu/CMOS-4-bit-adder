magic
tech scmos
timestamp 1578069705
<< nwell >>
rect -8 8 24 42
<< ntransistor >>
rect 3 -6 5 2
rect 11 -6 13 2
<< ptransistor >>
rect 3 14 5 34
rect 11 14 13 34
<< ndiffusion >>
rect 2 -6 3 2
rect 5 -6 11 2
rect 13 -6 14 2
<< pdiffusion >>
rect 2 14 3 34
rect 5 14 6 34
rect 10 14 11 34
rect 13 14 14 34
<< ndcontact >>
rect -2 -6 2 2
rect 14 -6 18 2
<< pdcontact >>
rect -2 14 2 34
rect 6 14 10 34
rect 14 14 18 34
<< polysilicon >>
rect 3 34 5 37
rect 11 34 13 37
rect 3 2 5 14
rect 11 2 13 14
rect 3 -9 5 -6
rect 11 -9 13 -6
<< metal1 >>
rect -8 38 24 42
rect -2 34 2 38
rect 14 34 18 38
rect 6 10 10 14
rect 6 6 24 10
rect 14 2 18 6
rect -2 -10 2 -6
rect -8 -14 24 -10
<< labels >>
rlabel metal1 0 39 0 39 5 vdd
rlabel metal1 4 -12 4 -12 1 gnd
rlabel polysilicon 4 36 4 36 1 a
rlabel polysilicon 12 36 12 36 1 b
rlabel metal1 22 8 22 8 7 out
<< end >>
